module top;
import uvm_pkg::*;
import tinyalu_pkg::*;
`include "uvm_macros.svh"
`include "tinyalu_pkg.svh"


endmodule : top